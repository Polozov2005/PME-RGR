.MODEL MBRM120L D(IS=1.52E-8 N=0.638 BV=20
+ IBV=0.0004 RS=0.0406 CJ=3E-10 VJ=0.374 MJ=0.379
+ TT=0.0)