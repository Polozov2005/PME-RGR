library IEEE;
use IEEE.std_logic_1164.all;

package mcu_functions is

  procedure  _pic_class( a: STD_LOGIC );
  procedure  _i8051_class( a: STD_LOGIC );
  procedure  _AVR_class( a: STD_LOGIC );
  procedure  _PIC18_class( a: STD_LOGIC );
  procedure  _MCP2515_class( a: STD_LOGIC );
  
end;

